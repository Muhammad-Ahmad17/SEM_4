library verilog;
use verilog.vl_types.all;
entity FSMdiv_vlg_vec_tst is
end FSMdiv_vlg_vec_tst;
