library verilog;
use verilog.vl_types.all;
entity FSM_sequence_detactor_vlg_vec_tst is
end FSM_sequence_detactor_vlg_vec_tst;
