LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

package My_Package is
	 component myDLatch is
		  port (
			clk   : in std_logic;
			D     : in std_logic;
			Q     : out std_logic;
			Q_not : out std_logic
			);
	end component;
end package My_Package;