library verilog;
use verilog.vl_types.all;
entity ahm_vlg_vec_tst is
end ahm_vlg_vec_tst;
