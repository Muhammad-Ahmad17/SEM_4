--------------SEVEN SEGMENT DISPLAY
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.my_compo.all;

entity fortuneWheel is 
	port (
        fpga_clk    : in  std_logic;
		  reset  : in std_logic;
        start_sw : in  std_logic;
		  led    : out std_logic_vector(7 downto 0);
        ssd0, ssd1, ssd2, ssd3 : out std_logic_vector(6 downto 0)
    );
end fortuneWheel;

architecture bhv of fortuneWheel is 
	--signals
   signal sclk, fclk : std_logic;
	signal ledout  : std_logic_vector(7 downto 0) := "00000001";
	signal ssdout  : std_logic_vector(6 downto 0) := "0000000";
	signal count   : std_logic_vector(31 downto 0) := X"00000000";
   signal input   : std_logic_vector(15 downto 0) := X"0000";  -- in hex  (fcount)
   --signal countSpeed : std_logic_vector(3 downto 0);
		
begin 
	---
	process (fpga_clk,start_sw)
	begin
		if (rising_edge(fpga_clk) and start_sw = '1') then 
		count <= count + 1;
		end if;
		fclk <= count(8);
		sclk <= count(22);
	end process;
	--- 
	
	--Slow Clock
    process (sclk,reset) is
    begin
			if reset = '1' then 
				ledout <=  "00000001";
			else
            ledout <= ledout(6 downto 0) & ledout(7);
        end if;
    end process;
	---	
	 --Fast Counter
    process (fclk,reset)
    begin
			if reset='1' then 
				input <= "0000000000000000";
        else
            input <= input + 1;
        end if;
    end process;
	 
	
	---
--	 u3: seven_seg port map (
--        bininput => input(15 downto 12),
--        cathodes => ssd3    
--    );
--    u2: seven_seg port map (
--        bininput => input(11 downto 8),
--        cathodes => ssd2    
--    );
--    u1: seven_seg port map (
--        bininput => input(7 downto 4),
--        cathodes => ssd1    
--    );
--    u0: seven_seg port map (
--        bininput => input(3 downto 0),
--        cathodes => ssd0    
--    );
process(input)
begin
    seven_seg(input(15 downto 12), ssd3);
    seven_seg(input(11 downto 8), ssd2);
    seven_seg(input(7 downto 4), ssd1);
    seven_seg(input(3 downto 0), ssd0);
end process;

	---
	led <= ledout;
end bhv;