library verilog;
use verilog.vl_types.all;
entity fortuneWheel_vlg_vec_tst is
end fortuneWheel_vlg_vec_tst;
