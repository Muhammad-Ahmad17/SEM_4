library verilog;
use verilog.vl_types.all;
entity ledBlinking_vlg_vec_tst is
end ledBlinking_vlg_vec_tst;
