library verilog;
use verilog.vl_types.all;
entity FSM_sequence_detactor_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FSM_sequence_detactor_vlg_check_tst;
